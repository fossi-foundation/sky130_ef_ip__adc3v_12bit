magic
tech sky130A
magscale 1 2
timestamp 1740521952
<< metal1 >>
rect 178772 36308 178936 36344
rect 176338 34661 178897 34697
<< metal2 >>
rect 175498 34596 175994 34978
rect 176423 34652 176523 35134
rect 177592 34816 177798 34962
rect 175492 34516 176029 34596
rect 173158 34315 173359 34488
rect 173564 34486 173664 34488
rect 173182 34204 173282 34315
rect 173517 34092 173718 34486
rect 173564 33962 173664 34092
rect 175492 32915 175555 34516
rect 175954 32915 176029 34516
rect 175492 32840 176029 32915
rect 176576 34528 177798 34816
rect 176576 32927 176639 34528
rect 177038 34500 177798 34528
rect 177038 32927 177113 34500
rect 176576 32835 177113 32927
rect 135656 7768 135691 8735
rect 138142 7892 138178 8738
rect 140678 8049 140706 8742
rect 143162 8179 143190 8762
rect 145650 8329 145678 8734
rect 148154 8455 148182 8756
rect 150644 8610 150672 8784
rect 153134 8621 153162 8740
rect 150644 8582 152284 8610
rect 148154 8427 152172 8455
rect 145650 8301 152060 8329
rect 143162 8151 151948 8179
rect 140678 8021 151836 8049
rect 138142 7856 150262 7892
rect 135656 7733 150079 7768
rect 150044 5987 150079 7733
rect 150043 5809 150079 5987
rect 150226 5802 150262 7856
rect 151808 5800 151836 8021
rect 151920 5800 151948 8151
rect 152032 5800 152060 8301
rect 152144 5800 152172 8427
rect 152256 5800 152284 8582
rect 152368 8593 153162 8621
rect 152368 5800 152396 8593
rect 155632 8462 155660 8760
rect 152480 8434 155660 8462
rect 152480 5800 152508 8434
rect 158136 8311 158164 8744
rect 152592 8283 158164 8311
rect 152592 5800 152620 8283
rect 160636 8173 160664 8748
rect 152704 8145 160664 8173
rect 152704 5800 152732 8145
rect 163126 8043 163154 8822
rect 152816 8015 163154 8043
rect 152816 5800 152844 8015
rect 165622 7900 165650 8750
rect 152928 7872 165650 7900
rect 152928 5800 152956 7872
rect 168122 7764 168150 8802
rect 153040 7736 168150 7764
rect 153040 5800 153068 7736
<< via2 >>
rect 172032 39160 172618 45534
rect 177978 34978 178524 45482
rect 175555 32915 175954 34516
rect 176639 32927 177038 34528
<< metal3 >>
rect 134771 61171 170336 61522
rect 134771 59799 135122 61171
rect 169985 60834 170336 61171
rect 169982 60815 170336 60834
rect 169982 59971 170005 60815
rect 170314 59971 170336 60815
rect 169982 59635 170336 59971
rect 169982 59284 170332 59635
rect 134422 48721 134588 48856
rect 171996 45534 172688 45626
rect 171996 39160 172032 45534
rect 172618 39160 172688 45534
rect 171996 39078 172688 39160
rect 177916 45482 178604 45570
rect 177916 34978 177978 45482
rect 178524 34978 178604 45482
rect 177916 34894 178604 34978
rect 175492 34516 176029 34596
rect 170234 34226 173282 34288
rect 170873 33979 173581 34041
rect 174067 33802 174129 34295
rect 170913 33778 174129 33802
rect 170913 33740 171728 33778
rect 171700 33678 171728 33740
rect 172692 33740 174129 33778
rect 172692 33678 172720 33740
rect 171700 33654 172720 33678
rect 175492 32915 175555 34516
rect 175954 32915 176029 34516
rect 175492 32840 176029 32915
rect 176576 34528 177113 34591
rect 176576 32927 176639 34528
rect 177038 32927 177113 34528
rect 176576 32835 177113 32927
<< via3 >>
rect 153572 60458 156089 60810
rect 149103 59834 151655 60183
rect 170005 59971 170314 60815
rect 152836 59432 153663 59589
rect 151777 59131 152604 59288
rect 172032 39160 172618 45534
rect 177978 34978 178524 45482
rect 171728 33678 172692 33778
rect 175555 32915 175954 34516
rect 176639 32927 177038 34528
rect 148574 10488 149640 10809
rect 156116 9884 157197 10215
<< metal4 >>
rect 149076 62401 151681 62578
rect 149076 61086 149206 62401
rect 151557 61086 151681 62401
rect 149076 60183 151681 61086
rect 149076 59834 149103 60183
rect 151655 59834 151681 60183
rect 149076 59795 151681 59834
rect 151934 59300 152385 64462
rect 152856 59600 153296 64473
rect 153550 64347 156115 64465
rect 153550 63032 153658 64347
rect 156009 63032 156115 64347
rect 153550 60810 156115 63032
rect 153550 60458 153572 60810
rect 156089 60458 156115 60810
rect 153550 60423 156115 60458
rect 169978 60815 170346 64471
rect 173564 64334 174584 64460
rect 173564 63007 173620 64334
rect 174483 63007 174584 64334
rect 169978 59971 170005 60815
rect 170314 59971 170346 60815
rect 169978 59949 170346 59971
rect 171701 62399 172721 62662
rect 171701 61072 171769 62399
rect 172632 61072 172721 62399
rect 152821 59589 153678 59600
rect 152821 59432 152836 59589
rect 153663 59432 153678 59589
rect 152821 59418 153678 59432
rect 151763 59288 152620 59300
rect 151763 59131 151777 59288
rect 152604 59131 152620 59288
rect 151763 59118 152620 59131
rect 134194 48721 134581 48856
rect 171701 45534 172721 61072
rect 173564 46879 174584 63007
rect 173564 46493 178605 46879
rect 173565 46116 178605 46493
rect 171701 39160 172032 45534
rect 172618 39160 172721 45534
rect 134194 35010 134447 35162
rect 171701 33802 172721 39160
rect 177842 45482 178605 46116
rect 177842 34978 177978 45482
rect 178524 34978 178605 45482
rect 177842 34873 178605 34978
rect 171700 33778 172721 33802
rect 171700 33678 171728 33778
rect 172692 33678 172721 33778
rect 171700 33654 172721 33678
rect 175492 34516 176029 34596
rect 175492 32915 175555 34516
rect 175954 32915 176029 34516
rect 175492 32779 176029 32915
rect 171701 32242 176029 32779
rect 176576 34528 177113 34591
rect 176576 32927 176639 34528
rect 177038 32927 177113 34528
rect 148524 10809 149674 10843
rect 148524 10488 148574 10809
rect 149640 10488 149674 10809
rect 148524 7274 149674 10488
rect 156059 10215 157241 10309
rect 156059 9884 156116 10215
rect 157197 9884 157241 10215
rect 156059 9849 157241 9884
rect 156076 9168 157235 9849
rect 156076 7817 156181 9168
rect 157121 7817 157235 9168
rect 156076 7713 157235 7817
rect 148524 5923 148622 7274
rect 149562 5923 149674 7274
rect 148524 5780 149674 5923
rect 171701 7340 172721 32242
rect 176576 31673 177113 32927
rect 173431 31136 177113 31673
rect 173431 9271 174450 31136
rect 173431 7799 173469 9271
rect 174416 7799 174450 9271
rect 173431 7725 174450 7799
rect 171701 5869 171750 7340
rect 172674 5869 172721 7340
rect 171701 5781 172721 5869
<< via4 >>
rect 149206 61086 151557 62401
rect 153658 63032 156009 64347
rect 173620 63007 174483 64334
rect 171769 61072 172632 62399
rect 156181 7817 157121 9168
rect 148622 5923 149562 7274
rect 173469 7799 174416 9271
rect 171750 5869 172674 7340
<< metal5 >>
rect 134194 64347 174641 64430
rect 134194 63032 153658 64347
rect 156009 64334 174641 64347
rect 156009 63032 173620 64334
rect 134194 63007 173620 63032
rect 174483 63007 174641 64334
rect 134194 62936 174641 63007
rect 134194 62401 174641 62495
rect 134194 61086 149206 62401
rect 151557 62399 174641 62401
rect 151557 61086 171769 62399
rect 134194 61072 171769 61086
rect 172632 61072 174641 62399
rect 134194 61001 174641 61072
rect 134194 9271 174457 9306
rect 134194 9168 173469 9271
rect 134194 7817 156181 9168
rect 157121 7817 173469 9168
rect 134194 7799 173469 7817
rect 174416 7799 174457 9271
rect 134194 7738 174457 7799
rect 134194 7340 174481 7381
rect 134194 7274 171750 7340
rect 134194 5923 148622 7274
rect 149562 5923 171750 7274
rect 134194 5869 171750 5923
rect 172674 5869 174481 7340
rect 134194 5813 174481 5869
use adc_via2_8cut  adc_via2_8cut_0
timestamp 1719106786
transform 0 -1 235996 1 0 27096
box 6850 62208 6998 62544
use adc_via2_8cut  adc_via2_8cut_1
timestamp 1719106786
transform 0 -1 235604 1 0 27336
box 6850 62208 6998 62544
use adc_via_3cut  adc_via_3cut_2
timestamp 1719452912
transform 0 1 69354 -1 0 45312
box 10601 106968 10663 107172
use sky130_ef_ip__cdac3v_12bit  sky130_ef_ip__cdac3v_12bit_0 ../ip/sky130_ef_ip__cdac3v_12bit/mag
timestamp 1731117925
transform 1 0 81345 0 -1 24388
box 52849 -36568 89580 15691
use sky130_ef_ip__scomp3v  sky130_ef_ip__scomp3v_0 ../ip/sky130_ef_ip__ccomp3v/mag
timestamp 1731034391
transform 0 1 174786 -1 0 45638
box -58 -3122 11186 4094
<< labels >>
flabel metal5 134965 61118 136829 62382 0 FreeSans 1600 0 0 0 vssa0
port 21 nsew ground bidirectional
flabel metal5 134951 63058 136815 64322 0 FreeSans 1600 0 0 0 vdda0
port 22 nsew power bidirectional
flabel metal1 178832 36308 178936 36344 0 FreeSans 320 180 0 0 adc0_ena
port 13 nsew signal input
flabel metal3 173139 34007 173148 34015 0 FreeSans 800 0 0 0 adc_aval
flabel metal1 178760 34661 178897 34697 0 FreeSans 320 180 0 0 adc0_comp_out
port 15 nsew signal output
flabel metal2 151808 5800 151836 6100 0 FreeSans 240 90 0 0 adc0_dac_val_0
port 12 nsew signal input
flabel metal2 151920 5800 151948 6100 0 FreeSans 240 90 0 0 adc0_dac_val_1
port 11 nsew signal input
flabel metal2 152032 5800 152060 6100 0 FreeSans 240 90 0 0 adc0_dac_val_2
port 10 nsew signal input
flabel metal2 152144 5800 152172 6100 0 FreeSans 240 90 0 0 adc0_dac_val_3
port 9 nsew signal input
flabel metal2 152256 5800 152284 6100 0 FreeSans 240 90 0 0 adc0_dac_val_4
port 8 nsew signal input
flabel metal2 152368 5800 152396 6100 0 FreeSans 240 90 0 0 adc0_dac_val_5
port 7 nsew signal input
flabel metal2 152480 5800 152508 6100 0 FreeSans 240 90 0 0 adc0_dac_val_6
port 6 nsew signal input
flabel metal2 152592 5800 152620 6100 0 FreeSans 240 90 0 0 adc0_dac_val_7
port 5 nsew signal input
flabel metal2 152704 5800 152732 6100 0 FreeSans 240 90 0 0 adc0_dac_val_8
port 4 nsew signal input
flabel metal2 152816 5800 152844 6100 0 FreeSans 240 90 0 0 adc0_dac_val_9
port 3 nsew signal input
flabel metal2 152928 5800 152956 6100 0 FreeSans 240 90 0 0 adc0_dac_val_10
port 2 nsew signal input
flabel metal2 153040 5800 153068 6100 0 FreeSans 240 90 0 0 adc0_dac_val_11
port 1 nsew signal input
flabel metal2 150043 5809 150079 5947 0 FreeSans 320 270 0 0 adc0_hold
port 16 nsew signal input
flabel metal2 150226 5802 150262 5956 0 FreeSans 320 90 0 0 adc0_reset
port 14 nsew signal input
flabel metal5 170392 7738 171538 9304 0 FreeSans 1600 0 0 0 vccd0
port 18 nsew power bidirectional
flabel metal5 170486 5813 171529 7379 0 FreeSans 1600 0 0 0 vssd0
port 19 nsew ground bidirectional
flabel metal4 151953 64262 152328 64462 0 FreeSans 320 0 0 0 adc_vrefL
port 17 nsew analog bidirectional
flabel metal4 152925 64273 153181 64473 0 FreeSans 320 0 0 0 adc_vrefH
port 20 nsew analog bidirectional
flabel metal4 169978 63893 170345 64471 0 FreeSans 1600 0 0 0 adc_vCM
port 24 nsew analog bidirectional
flabel metal4 134194 48721 134360 48856 0 FreeSans 1600 0 0 0 adc_trim
port 23 nsew analog input
flabel metal4 134194 35010 134447 35162 0 FreeSans 1600 0 0 0 adc0
port 25 nsew analog input
<< end >>
