magic
tech sky130A
magscale 1 2
timestamp 1740586040
<< metal2 >>
rect 41304 28796 41800 29178
rect 42229 28852 42329 29334
rect 43398 29016 43604 29162
rect 41298 28716 41835 28796
rect 38964 28515 39165 28688
rect 39370 28686 39470 28688
rect 38988 28404 39088 28515
rect 39323 28292 39524 28686
rect 39370 28162 39470 28292
rect 41298 27115 41361 28716
rect 41760 27115 41835 28716
rect 41298 27040 41835 27115
rect 42382 28728 43604 29016
rect 42382 27127 42445 28728
rect 42844 28700 43604 28728
rect 42844 27127 42919 28700
rect 42382 27035 42919 27127
rect 1462 1968 1497 2935
rect 3948 2092 3984 2938
rect 6484 2249 6512 2942
rect 8968 2379 8996 2962
rect 11456 2529 11484 2934
rect 13960 2655 13988 2956
rect 16450 2810 16478 2984
rect 18940 2821 18968 2940
rect 16450 2782 18090 2810
rect 13960 2627 17978 2655
rect 11456 2501 17866 2529
rect 8968 2351 17754 2379
rect 6484 2221 17642 2249
rect 3948 2056 16068 2092
rect 1462 1933 15885 1968
rect 15850 187 15885 1933
rect 15849 0 15885 187
rect 16032 0 16068 2056
rect 17614 0 17642 2221
rect 17726 0 17754 2351
rect 17838 0 17866 2501
rect 17950 0 17978 2627
rect 18062 0 18090 2782
rect 18174 2793 18968 2821
rect 18174 0 18202 2793
rect 21438 2662 21466 2960
rect 18286 2634 21466 2662
rect 18286 0 18314 2634
rect 23942 2511 23970 2944
rect 18398 2483 23970 2511
rect 18398 0 18426 2483
rect 26442 2373 26470 2948
rect 18510 2345 26470 2373
rect 18510 0 18538 2345
rect 28932 2243 28960 3022
rect 18622 2215 28960 2243
rect 18622 0 18650 2215
rect 31428 2100 31456 2950
rect 18734 2072 31456 2100
rect 18734 0 18762 2072
rect 33928 1964 33956 3002
rect 18846 1936 33956 1964
rect 18846 0 18874 1936
<< via2 >>
rect 37838 33360 38424 39734
rect 43784 29178 44330 39682
rect 41361 27115 41760 28716
rect 42445 27127 42844 28728
<< metal3 >>
rect 577 55371 36142 55722
rect 577 53999 928 55371
rect 35791 55034 36142 55371
rect 35788 55015 36142 55034
rect 35788 54171 35811 55015
rect 36120 54171 36142 55015
rect 35788 53835 36142 54171
rect 35788 53484 36138 53835
rect 0 42921 394 43056
rect 37802 39734 38494 39826
rect 37802 33360 37838 39734
rect 38424 33360 38494 39734
rect 37802 33278 38494 33360
rect 43722 39682 44410 39770
rect 0 29210 259 29362
rect 43722 29178 43784 39682
rect 44330 29178 44410 39682
rect 44578 30496 44742 30558
rect 43722 29094 44410 29178
rect 42144 28861 44703 28921
rect 41298 28716 41835 28796
rect 36040 28426 39088 28488
rect 36679 28179 39387 28241
rect 39873 28002 39935 28495
rect 36719 27978 39935 28002
rect 36719 27940 37534 27978
rect 37506 27878 37534 27940
rect 38498 27940 39935 27978
rect 38498 27878 38526 27940
rect 37506 27854 38526 27878
rect 41298 27115 41361 28716
rect 41760 27115 41835 28716
rect 41298 27040 41835 27115
rect 42382 28728 42919 28791
rect 42382 27127 42445 28728
rect 42844 27127 42919 28728
rect 42382 27035 42919 27127
<< via3 >>
rect 19378 54658 21895 55010
rect 14909 54034 17461 54383
rect 35811 54171 36120 55015
rect 18642 53632 19469 53789
rect 17583 53331 18410 53488
rect 37838 33360 38424 39734
rect 43784 29178 44330 39682
rect 37534 27878 38498 27978
rect 41361 27115 41760 28716
rect 42445 27127 42844 28728
rect 14380 4688 15446 5009
rect 21922 4084 23003 4415
<< metal4 >>
rect 14882 56601 17487 56778
rect 14882 55286 15012 56601
rect 17363 55286 17487 56601
rect 14882 54383 17487 55286
rect 14882 54034 14909 54383
rect 17461 54034 17487 54383
rect 14882 53995 17487 54034
rect 17740 53500 18191 58662
rect 18651 53800 19102 58673
rect 19356 58547 21921 58665
rect 19356 57232 19464 58547
rect 21815 57232 21921 58547
rect 19356 55010 21921 57232
rect 19356 54658 19378 55010
rect 21895 54658 21921 55010
rect 19356 54623 21921 54658
rect 35784 55015 36152 58671
rect 39370 58534 40390 58660
rect 39370 57207 39426 58534
rect 40289 57207 40390 58534
rect 35784 54171 35811 55015
rect 36120 54171 36152 55015
rect 35784 54149 36152 54171
rect 37507 56599 38527 56862
rect 37507 55272 37575 56599
rect 38438 55272 38527 56599
rect 18627 53789 19484 53800
rect 18627 53632 18642 53789
rect 19469 53632 19484 53789
rect 18627 53618 19484 53632
rect 17569 53488 18426 53500
rect 17569 53331 17583 53488
rect 18410 53331 18426 53488
rect 17569 53318 18426 53331
rect 37507 39734 38527 55272
rect 39370 41079 40390 57207
rect 39370 40693 44411 41079
rect 39371 40316 44411 40693
rect 37507 33360 37838 39734
rect 38424 33360 38527 39734
rect 37507 28002 38527 33360
rect 43648 39682 44411 40316
rect 43648 29178 43784 39682
rect 44330 29178 44411 39682
rect 43648 29073 44411 29178
rect 37506 27978 38527 28002
rect 37506 27878 37534 27978
rect 38498 27878 38527 27978
rect 37506 27854 38527 27878
rect 41298 28716 41835 28796
rect 41298 27115 41361 28716
rect 41760 27115 41835 28716
rect 41298 26979 41835 27115
rect 37507 26442 41835 26979
rect 42382 28728 42919 28791
rect 42382 27127 42445 28728
rect 42844 27127 42919 28728
rect 14330 5009 15480 5043
rect 14330 4688 14380 5009
rect 15446 4688 15480 5009
rect 14330 1474 15480 4688
rect 21865 4415 23047 4509
rect 21865 4084 21922 4415
rect 23003 4084 23047 4415
rect 21865 4049 23047 4084
rect 21882 3368 23041 4049
rect 21882 2017 21987 3368
rect 22927 2017 23041 3368
rect 21882 1913 23041 2017
rect 14330 123 14428 1474
rect 15368 123 15480 1474
rect 14330 13 15480 123
rect 37507 1540 38527 26442
rect 42382 25873 42919 27127
rect 39237 25336 42919 25873
rect 39237 3471 40256 25336
rect 39237 1999 39275 3471
rect 40222 1999 40256 3471
rect 39237 1938 40256 1999
rect 37507 69 37556 1540
rect 38480 69 38527 1540
rect 37507 13 38527 69
<< via4 >>
rect 15012 55286 17363 56601
rect 19464 57232 21815 58547
rect 39426 57207 40289 58534
rect 37575 55272 38438 56599
rect 21987 2017 22927 3368
rect 14428 123 15368 1474
rect 39275 1999 40222 3471
rect 37556 69 38480 1540
<< metal5 >>
rect 0 58547 40447 58630
rect 0 57232 19464 58547
rect 21815 58534 40447 58547
rect 21815 57232 39426 58534
rect 0 57207 39426 57232
rect 40289 57207 40447 58534
rect 0 57136 40447 57207
rect 0 56601 40447 56695
rect 0 55286 15012 56601
rect 17363 56599 40447 56601
rect 17363 55286 37575 56599
rect 0 55272 37575 55286
rect 38438 55272 40447 56599
rect 0 55201 40447 55272
rect 0 3471 40263 3506
rect 0 3368 39275 3471
rect 0 2017 21987 3368
rect 22927 2017 39275 3368
rect 0 1999 39275 2017
rect 40222 1999 40263 3471
rect 0 1938 40263 1999
rect 0 1540 40287 1581
rect 0 1474 37556 1540
rect 0 123 14428 1474
rect 15368 123 37556 1474
rect 0 69 37556 123
rect 38480 69 40287 1540
rect 0 13 40287 69
use adc_via2_8cut  adc_via2_8cut_0
timestamp 1719106786
transform 0 -1 101802 1 0 21296
box 6850 62208 6998 62544
use adc_via2_8cut  adc_via2_8cut_1
timestamp 1719106786
transform 0 -1 101410 1 0 21536
box 6850 62208 6998 62544
use adc_via2_8cut  adc_via2_8cut_2
timestamp 1719106786
transform -1 0 51490 0 -1 92905
box 6850 62208 6998 62544
use adc_via2_8cut  adc_via2_8cut_3
timestamp 1719106786
transform 0 1 -20216 -1 0 35840
box 6850 62208 6998 62544
use adc_via_3cut  adc_via_3cut_2
timestamp 1719452912
transform -1 0 55203 0 -1 137594
box 10601 106968 10663 107172
use sky130_ef_ip__cdac3v_12bit  sky130_ef_ip__cdac3v_12bit_0 ../ip/sky130_ef_ip__cdac3v_12bit/mag
timestamp 1731117925
transform 1 0 -52849 0 -1 18588
box 52849 -36568 89580 15691
use sky130_ef_ip__scomp3v  sky130_ef_ip__scomp3v_0 ../ip/sky130_ef_ip__ccomp3v/mag
timestamp 1731034391
transform 0 1 40592 -1 0 39838
box -58 -3122 11186 4094
<< labels >>
flabel metal5 s 0 55201 40447 56695 0 FreeSans 1600 0 0 0 vssa0
port 21 nsew ground bidirectional
flabel metal5 s 0 57136 40447 58630 0 FreeSans 1600 0 0 0 vdda0
port 22 nsew power bidirectional
flabel metal3 44616 30496 44742 30558 0 FreeSans 320 180 0 0 adc0_ena
port 13 nsew signal input
flabel metal3 38945 28207 38954 28215 0 FreeSans 800 0 0 0 adc_aval
flabel metal3 44566 28861 44703 28921 0 FreeSans 320 180 0 0 adc0_comp_out
port 15 nsew signal output
flabel metal2 17614 0 17642 300 0 FreeSans 240 90 0 0 adc0_dac_val_0
port 12 nsew signal input
flabel metal2 17726 0 17754 300 0 FreeSans 240 90 0 0 adc0_dac_val_1
port 11 nsew signal input
flabel metal2 17838 0 17866 300 0 FreeSans 240 90 0 0 adc0_dac_val_2
port 10 nsew signal input
flabel metal2 17950 0 17978 300 0 FreeSans 240 90 0 0 adc0_dac_val_3
port 9 nsew signal input
flabel metal2 18062 0 18090 300 0 FreeSans 240 90 0 0 adc0_dac_val_4
port 8 nsew signal input
flabel metal2 18174 0 18202 300 0 FreeSans 240 90 0 0 adc0_dac_val_5
port 7 nsew signal input
flabel metal2 18286 0 18314 300 0 FreeSans 240 90 0 0 adc0_dac_val_6
port 6 nsew signal input
flabel metal2 18398 0 18426 300 0 FreeSans 240 90 0 0 adc0_dac_val_7
port 5 nsew signal input
flabel metal2 18510 0 18538 300 0 FreeSans 240 90 0 0 adc0_dac_val_8
port 4 nsew signal input
flabel metal2 18622 0 18650 300 0 FreeSans 240 90 0 0 adc0_dac_val_9
port 3 nsew signal input
flabel metal2 18734 0 18762 300 0 FreeSans 240 90 0 0 adc0_dac_val_10
port 2 nsew signal input
flabel metal2 18846 0 18874 300 0 FreeSans 240 90 0 0 adc0_dac_val_11
port 1 nsew signal input
flabel metal2 15849 0 15885 300 0 FreeSans 320 270 0 0 adc0_hold
port 16 nsew signal input
flabel metal2 16032 0 16068 300 0 FreeSans 320 90 0 0 adc0_reset
port 14 nsew signal input
flabel metal5 s 0 1938 40263 3506 0 FreeSans 1600 0 0 0 vccd0
port 18 nsew power bidirectional
flabel metal5 s 0 13 40287 1581 0 FreeSans 1600 0 0 0 vssd0
port 19 nsew ground bidirectional
flabel metal4 17740 58047 18191 58662 0 FreeSans 320 0 0 0 adc_vrefL
port 17 nsew analog bidirectional
flabel metal4 18651 58058 19102 58673 0 FreeSans 320 0 0 0 adc_vrefH
port 20 nsew analog bidirectional
flabel metal4 35784 58093 36151 58671 0 FreeSans 1600 0 0 0 adc_vCM
port 24 nsew analog bidirectional
flabel metal3 0 29210 253 29362 0 FreeSans 1600 0 0 0 adc0
port 25 nsew analog input
flabel metal3 0 42921 166 43056 0 FreeSans 1600 0 0 0 adc_trim
port 23 nsew analog input
<< end >>
