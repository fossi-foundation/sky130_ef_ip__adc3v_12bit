VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__adc3v_12bit
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__adc3v_12bit ;
  ORIGIN -670.970 -28.900 ;
  SIZE 223.710 BY 293.465 ;
  PIN adc0_dac_val_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 765.200 29.000 765.340 38.820 ;
    END
  END adc0_dac_val_11
  PIN adc0_dac_val_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 764.640 29.000 764.780 39.500 ;
    END
  END adc0_dac_val_10
  PIN adc0_dac_val_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 764.080 29.000 764.220 40.215 ;
    END
  END adc0_dac_val_9
  PIN adc0_dac_val_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 763.520 29.000 763.660 40.865 ;
    END
  END adc0_dac_val_8
  PIN adc0_dac_val_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 762.960 29.000 763.100 41.555 ;
    END
  END adc0_dac_val_7
  PIN adc0_dac_val_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 762.400 29.000 762.540 42.310 ;
    END
  END adc0_dac_val_6
  PIN adc0_dac_val_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 761.840 29.000 761.980 43.105 ;
    END
  END adc0_dac_val_5
  PIN adc0_dac_val_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 761.280 29.000 761.420 43.050 ;
    END
  END adc0_dac_val_4
  PIN adc0_dac_val_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 760.720 29.000 760.860 42.275 ;
    END
  END adc0_dac_val_3
  PIN adc0_dac_val_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 760.160 29.000 760.300 41.645 ;
    END
  END adc0_dac_val_2
  PIN adc0_dac_val_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 759.600 29.000 759.740 40.895 ;
    END
  END adc0_dac_val_1
  PIN adc0_dac_val_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 759.040 29.000 759.180 40.245 ;
    END
  END adc0_dac_val_0
  PIN adc0_ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met1 ;
        RECT 891.675 181.540 894.680 181.720 ;
    END
  END adc0_ena
  PIN adc0_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 751.130 29.010 751.310 39.460 ;
    END
  END adc0_reset
  PIN adc0_comp_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met1 ;
        RECT 882.600 173.305 894.485 173.485 ;
    END
  END adc0_comp_out
  PIN adc0_hold
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 750.215 29.045 750.395 29.935 ;
    END
  END adc0_hold
  PIN adc_vrefL
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 121.799995 ;
    PORT
      LAYER met4 ;
        RECT 759.670 296.440 761.925 322.310 ;
    END
  END adc_vrefL
  PIN vccd0
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 785.605 38.690 867.345 46.530 ;
    END
  END vccd0
  PIN vssd0
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 747.810 29.065 858.750 36.905 ;
    END
  END vssd0
  PIN adc_vrefH
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 121.799995 ;
    PORT
      LAYER met4 ;
        RECT 764.280 297.945 766.480 322.365 ;
    END
  END adc_vrefH
  PIN vssa0
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 670.970 305.005 746.030 312.475 ;
    END
  END vssa0
  PIN vdda0
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 670.970 314.680 768.290 322.150 ;
    END
  END vdda0
  PIN adc_trim
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 670.970 243.605 672.940 244.280 ;
    END
  END adc_trim
  PIN adc_vCM
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNAGATEAREA 70.000000 ;
    ANTENNADIFFAREA 121.799995 ;
    PORT
      LAYER met4 ;
        RECT 849.890 304.075 851.730 322.355 ;
    END
  END adc_vCM
  PIN adc0
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 10.440000 ;
    PORT
      LAYER met4 ;
        RECT 670.970 175.050 672.265 175.810 ;
    END
  END adc0
  OBS
      LAYER nwell ;
        RECT 673.165 43.775 894.400 295.200 ;
      LAYER li1 ;
        RECT 673.600 43.905 894.070 294.810 ;
      LAYER met1 ;
        RECT 670.970 182.000 894.070 298.945 ;
        RECT 670.970 181.260 891.395 182.000 ;
        RECT 670.970 173.765 894.070 181.260 ;
        RECT 670.970 173.025 882.320 173.765 ;
        RECT 670.970 43.875 894.070 173.025 ;
      LAYER met2 ;
        RECT 671.005 43.385 892.860 304.780 ;
        RECT 671.005 43.330 761.560 43.385 ;
        RECT 671.005 42.555 761.000 43.330 ;
        RECT 762.260 42.590 892.860 43.385 ;
        RECT 671.005 41.925 760.440 42.555 ;
        RECT 671.005 41.175 759.880 41.925 ;
        RECT 762.820 41.835 892.860 42.590 ;
        RECT 671.005 40.525 759.320 41.175 ;
        RECT 763.380 41.145 892.860 41.835 ;
        RECT 671.005 39.740 758.760 40.525 ;
        RECT 763.940 40.495 892.860 41.145 ;
        RECT 764.500 39.780 892.860 40.495 ;
        RECT 671.005 30.215 750.850 39.740 ;
        RECT 671.005 29.935 749.935 30.215 ;
        RECT 750.675 29.935 750.850 30.215 ;
        RECT 751.590 29.935 758.760 39.740 ;
        RECT 765.060 39.100 892.860 39.780 ;
        RECT 765.620 29.935 892.860 39.100 ;
      LAYER met3 ;
        RECT 672.110 47.230 893.020 307.610 ;
      LAYER met4 ;
        RECT 672.205 296.040 759.270 322.325 ;
        RECT 762.325 297.545 763.880 322.325 ;
        RECT 766.880 303.675 849.490 322.325 ;
        RECT 852.130 303.675 893.025 322.325 ;
        RECT 766.880 297.545 893.025 303.675 ;
        RECT 762.325 296.040 893.025 297.545 ;
        RECT 672.205 244.680 893.025 296.040 ;
        RECT 673.340 243.205 893.025 244.680 ;
        RECT 672.205 176.210 893.025 243.205 ;
        RECT 672.665 174.650 893.025 176.210 ;
        RECT 672.205 28.900 893.025 174.650 ;
      LAYER met5 ;
        RECT 769.890 313.080 873.205 322.150 ;
        RECT 747.630 303.405 873.205 313.080 ;
        RECT 670.970 48.130 873.205 303.405 ;
        RECT 670.970 46.530 784.005 48.130 ;
        RECT 670.970 45.840 785.605 46.530 ;
        RECT 670.970 39.085 784.005 45.840 ;
        RECT 670.970 38.690 785.605 39.085 ;
        RECT 670.970 38.505 784.005 38.690 ;
        RECT 670.970 36.905 746.210 38.505 ;
        RECT 868.945 37.090 873.205 48.130 ;
        RECT 670.970 36.370 747.810 36.905 ;
        RECT 670.970 29.615 746.210 36.370 ;
        RECT 670.970 29.065 747.810 29.615 ;
        RECT 860.350 29.065 873.205 37.090 ;
  END
END sky130_ef_ip__adc3v_12bit
END LIBRARY

