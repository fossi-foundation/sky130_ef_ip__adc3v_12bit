VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__adc3v_12bit
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__adc3v_12bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.710 BY 293.365 ;
  PIN adc_dac_val[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 94.230 0.000 94.370 1.500 ;
    END
  END adc_dac_val[11]
  PIN adc_dac_val[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 93.670 0.000 93.810 1.500 ;
    END
  END adc_dac_val[10]
  PIN adc_dac_val[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 93.110 0.000 93.250 1.500 ;
    END
  END adc_dac_val[9]
  PIN adc_dac_val[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.690 1.500 ;
    END
  END adc_dac_val[8]
  PIN adc_dac_val[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 91.990 0.000 92.130 1.500 ;
    END
  END adc_dac_val[7]
  PIN adc_dac_val[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 91.430 0.000 91.570 1.500 ;
    END
  END adc_dac_val[6]
  PIN adc_dac_val[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 90.870 0.000 91.010 1.500 ;
    END
  END adc_dac_val[5]
  PIN adc_dac_val[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 90.310 0.000 90.450 1.500 ;
    END
  END adc_dac_val[4]
  PIN adc_dac_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 89.750 0.000 89.890 1.500 ;
    END
  END adc_dac_val[3]
  PIN adc_dac_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 89.190 0.000 89.330 1.500 ;
    END
  END adc_dac_val[2]
  PIN adc_dac_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 88.630 0.000 88.770 1.500 ;
    END
  END adc_dac_val[1]
  PIN adc_dac_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 88.070 0.000 88.210 1.500 ;
    END
  END adc_dac_val[0]
  PIN adc_ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met1 ;
        RECT 222.700 152.375 223.010 153.130 ;
        RECT 222.570 152.010 223.570 152.375 ;
        RECT 222.210 151.750 223.570 152.010 ;
        RECT 222.570 151.375 223.570 151.750 ;
      LAYER met2 ;
        RECT 222.460 151.805 223.200 153.485 ;
      LAYER met3 ;
        RECT 222.460 152.790 223.200 153.485 ;
        RECT 222.460 152.480 223.710 152.790 ;
        RECT 222.460 151.805 223.200 152.480 ;
    END
  END adc_ena
  PIN adc_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 80.160 0.000 80.340 1.500 ;
    END
  END adc_reset
  PIN adc_comp_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met3 ;
        RECT 222.210 144.305 223.515 144.605 ;
    END
  END adc_comp_out
  PIN adc_hold
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.859200 ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER met2 ;
        RECT 79.245 0.000 79.425 1.500 ;
    END
  END adc_hold
  PIN adc_vrefL
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 121.799995 ;
    PORT
      LAYER met4 ;
        RECT 88.700 290.235 90.955 293.310 ;
    END
  END adc_vrefL
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 71.650 0.065 77.400 1.500 ;
        RECT 187.535 0.065 192.635 1.500 ;
      LAYER met5 ;
        RECT 0.000 0.065 201.435 7.905 ;
    END
  END vssd
  PIN adc_vrefH
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 121.799995 ;
    PORT
      LAYER met4 ;
        RECT 93.255 290.290 95.510 293.365 ;
    END
  END adc_vrefH
  PIN adc_trim
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.605 1.500 215.280 ;
    END
  END adc_trim
  PIN adc_vCM
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNAGATEAREA 70.000000 ;
    ANTENNADIFFAREA 121.799995 ;
    PORT
      LAYER met4 ;
        RECT 178.920 291.865 180.760 293.355 ;
        RECT 178.920 290.465 180.755 291.865 ;
    END
  END adc_vCM
  PIN adc_in
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 10.440000 ;
    PORT
      LAYER met3 ;
        RECT 1.235 146.810 1.500 148.805 ;
        RECT 0.000 146.050 1.500 146.810 ;
        RECT 1.235 144.750 1.500 146.050 ;
      LAYER met4 ;
        RECT 1.235 144.750 1.500 146.910 ;
    END
  END adc_in
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 9.690 201.315 17.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.185 9.690 201.280 129.365 ;
    END
  END vccd
  PIN vdda
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 222.210 155.820 223.670 199.720 ;
      LAYER li1 ;
        RECT 222.210 199.010 223.340 199.385 ;
        RECT 222.965 156.595 223.340 199.010 ;
        RECT 222.210 156.220 223.340 156.595 ;
      LAYER met1 ;
        RECT 222.210 199.010 223.340 199.385 ;
        RECT 222.965 156.595 223.340 199.010 ;
        RECT 222.210 156.220 223.340 156.595 ;
      LAYER met4 ;
        RECT 96.780 291.865 109.605 293.325 ;
        RECT 196.850 291.865 201.950 293.300 ;
      LAYER met5 ;
        RECT 0.000 285.680 202.235 293.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.240 145.365 222.055 205.395 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.950 201.580 218.240 205.395 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 276.005 202.235 283.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 187.530 139.270 192.635 284.310 ;
    END
  END vssa
  OBS
      LAYER nwell ;
        RECT 2.195 14.775 222.210 266.200 ;
      LAYER li1 ;
        RECT 2.630 14.905 222.210 265.810 ;
      LAYER met1 ;
        RECT 1.500 241.600 222.210 269.945 ;
        RECT 1.200 241.300 222.210 241.600 ;
        RECT 1.500 205.570 222.210 241.300 ;
        RECT 1.200 205.330 222.210 205.570 ;
        RECT 1.500 169.815 222.210 205.330 ;
        RECT 1.480 169.555 222.210 169.815 ;
        RECT 1.200 169.315 222.210 169.555 ;
        RECT 1.480 168.760 222.210 169.315 ;
        RECT 0.995 111.515 1.255 111.535 ;
        RECT 1.500 111.515 222.210 168.760 ;
        RECT 0.995 111.275 222.210 111.515 ;
        RECT 0.995 110.480 1.255 111.275 ;
        RECT 0.515 75.490 0.775 75.510 ;
        RECT 1.500 75.490 222.210 111.275 ;
        RECT 0.515 75.250 222.210 75.490 ;
        RECT 0.515 74.455 0.775 75.250 ;
        RECT 0.035 39.470 0.295 39.485 ;
        RECT 1.500 39.470 222.210 75.250 ;
        RECT 0.035 39.230 222.210 39.470 ;
        RECT 0.035 38.430 0.295 39.230 ;
        RECT 0.035 26.995 0.295 27.010 ;
        RECT 1.500 26.995 222.210 39.230 ;
        RECT 0.000 26.755 222.210 26.995 ;
        RECT 0.035 25.955 0.295 26.755 ;
        RECT 0.520 26.515 0.780 26.525 ;
        RECT 1.500 26.515 222.210 26.755 ;
        RECT 0.500 26.275 222.210 26.515 ;
        RECT 0.520 25.470 0.780 26.275 ;
        RECT 0.995 26.035 1.255 26.045 ;
        RECT 1.500 26.035 222.210 26.275 ;
        RECT 0.985 25.795 222.210 26.035 ;
        RECT 0.995 24.990 1.255 25.795 ;
        RECT 1.500 25.565 222.210 25.795 ;
        RECT 1.475 25.555 222.210 25.565 ;
        RECT 1.465 25.315 222.210 25.555 ;
        RECT 1.475 24.510 222.210 25.315 ;
        RECT 1.500 14.875 222.210 24.510 ;
      LAYER met2 ;
        RECT 1.500 169.815 222.130 275.780 ;
        RECT 1.480 168.760 222.130 169.815 ;
        RECT 0.995 110.480 1.255 111.535 ;
        RECT 0.530 75.510 0.770 75.515 ;
        RECT 0.515 74.455 0.775 75.510 ;
        RECT 0.050 39.485 0.290 39.490 ;
        RECT 0.035 38.430 0.295 39.485 ;
        RECT 0.050 27.010 0.290 38.430 ;
        RECT 0.035 25.955 0.295 27.010 ;
        RECT 0.530 26.525 0.770 74.455 ;
        RECT 0.520 25.470 0.780 26.525 ;
        RECT 1.010 26.045 1.250 110.480 ;
        RECT 0.995 24.990 1.255 26.045 ;
        RECT 1.490 25.565 222.130 168.760 ;
        RECT 1.475 24.510 222.130 25.565 ;
        RECT 1.500 1.500 222.130 24.510 ;
      LAYER met3 ;
        RECT 1.500 18.230 222.210 278.610 ;
      LAYER met4 ;
        RECT 1.500 1.500 214.595 291.865 ;
      LAYER met5 ;
        RECT 29.155 28.510 154.505 265.525 ;
  END
END sky130_ef_ip__adc3v_12bit
END LIBRARY

