magic
tech sky130A
timestamp 1719106786
<< checkpaint >>
rect 3425 31104 3499 31272
<< metal2 >>
rect 3425 31266 3499 31272
rect 3425 31110 3428 31266
rect 3496 31110 3499 31266
rect 3425 31104 3499 31110
<< via2 >>
rect 3428 31110 3496 31266
<< metal3 >>
rect 3425 31266 3499 31272
rect 3425 31110 3428 31266
rect 3496 31110 3499 31266
rect 3425 31104 3499 31110
<< end >>
