magic
tech sky130A
magscale 1 2
timestamp 1719173267
<< checkpaint >>
rect 566656 91154 566956 91980
<< metal3 >>
rect 566656 91972 566956 91980
rect 566656 91165 566665 91972
rect 566947 91165 566956 91972
rect 566656 91154 566956 91165
<< via3 >>
rect 566665 91165 566947 91972
<< metal4 >>
rect 566656 91972 566956 91980
rect 566656 91165 566665 91972
rect 566947 91165 566956 91972
rect 566656 91154 566956 91165
<< end >>
