magic
tech sky130A
magscale 1 2
timestamp 1719452912
<< checkpaint >>
rect 10601 106968 10663 107172
<< metal1 >>
rect 10601 107166 10663 107172
rect 10601 106974 10606 107166
rect 10658 106974 10663 107166
rect 10601 106968 10663 106974
<< via1 >>
rect 10606 106974 10658 107166
<< metal2 >>
rect 10601 107166 10663 107172
rect 10601 106974 10606 107166
rect 10658 106974 10663 107166
rect 10601 106968 10663 106974
<< end >>
