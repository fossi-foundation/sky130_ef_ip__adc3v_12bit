magic
tech sky130A
magscale 1 2
timestamp 1731119720
<< error_s >>
rect 167137 7822 167138 8242
rect 167197 7882 167198 8182
<< metal1 >>
rect 173946 28794 173952 28846
rect 174004 28838 174010 28846
rect 178204 28838 178240 28888
rect 174004 28802 178240 28838
rect 174004 28794 174010 28802
rect 135641 8585 135647 8637
rect 135699 8628 135705 8637
rect 173600 8628 173606 8636
rect 135699 8593 173606 8628
rect 135699 8585 135705 8593
rect 173600 8584 173606 8593
rect 173658 8584 173664 8636
rect 173946 8514 173952 8522
rect 136762 8478 173952 8514
rect 173946 8470 173952 8478
rect 174004 8470 174010 8522
rect 170288 1996 176422 2005
rect 170288 1969 176329 1996
rect 176381 1969 176422 1996
rect 173600 1921 173606 1928
rect 170288 1885 173606 1921
rect 173600 1876 173606 1885
rect 173658 1876 173664 1928
<< via1 >>
rect 173952 28794 174004 28846
rect 135647 8585 135699 8637
rect 173606 8584 173658 8636
rect 173952 8470 174004 8522
rect 173606 1876 173658 1928
<< metal2 >>
rect 175652 34288 176450 34388
rect 175678 33906 176510 34006
rect 175530 31718 176854 32100
rect 175530 31170 175911 31718
rect 173952 28846 174004 28852
rect 173952 28788 174004 28794
rect 135656 8643 135691 8735
rect 135647 8637 135699 8643
rect 135647 8579 135699 8585
rect 138142 6812 138178 8738
rect 140678 6969 140706 8742
rect 143162 7149 143190 8762
rect 145650 7299 145678 8734
rect 148154 7425 148182 8756
rect 150644 7580 150672 8784
rect 153134 8371 153162 8740
rect 152368 8343 153162 8371
rect 150644 7552 152284 7580
rect 148154 7397 152172 7425
rect 145650 7271 152060 7299
rect 143162 7121 151948 7149
rect 140678 6941 151836 6969
rect 138142 6776 150262 6812
rect 150226 102 150262 6776
rect 151808 0 151836 6941
rect 151920 0 151948 7121
rect 152032 0 152060 7271
rect 152144 0 152172 7397
rect 152256 0 152284 7552
rect 152368 0 152396 8343
rect 155632 8212 155660 8760
rect 152480 8184 155660 8212
rect 152480 0 152508 8184
rect 158136 8031 158164 8744
rect 152592 8003 158164 8031
rect 152592 0 152620 8003
rect 160636 7893 160664 8748
rect 152704 7865 160664 7893
rect 152704 0 152732 7865
rect 163126 7713 163154 8822
rect 152816 7685 163154 7713
rect 152816 0 152844 7685
rect 165622 7570 165650 8750
rect 152928 7542 165650 7570
rect 152928 0 152956 7542
rect 168122 7384 168150 8802
rect 173606 8636 173658 8642
rect 173606 8578 173658 8584
rect 153040 7356 168150 7384
rect 153040 0 153068 7356
rect 173614 1934 173649 8578
rect 173960 8528 173996 28788
rect 175529 27072 175911 31170
rect 176303 31060 176908 31160
rect 175498 26596 175994 27072
rect 175492 26516 176029 26596
rect 175492 24915 175555 26516
rect 175954 24915 176029 26516
rect 175492 24840 176029 24915
rect 173952 8522 174004 8528
rect 173952 8464 174004 8470
rect 176303 1996 176403 31060
rect 176528 29802 176848 30008
rect 176528 27308 176734 29802
rect 176528 26591 177082 27308
rect 176528 26528 177113 26591
rect 176528 26487 176639 26528
rect 176576 24927 176639 26487
rect 177038 24927 177113 26528
rect 176576 24835 177113 24927
rect 173606 1928 173658 1934
rect 173606 1870 173658 1876
rect 173614 1865 173649 1870
rect 176303 1804 176329 1996
rect 176381 1804 176403 1996
rect 176303 1794 176403 1804
<< via2 >>
rect 181062 34968 187436 35554
rect 175555 24915 175954 26516
rect 176910 29110 187414 29656
rect 176639 24927 177038 26528
<< metal3 >>
rect 180980 35554 187528 35590
rect 180980 34968 181062 35554
rect 187436 34968 187528 35554
rect 180980 34898 187528 34968
rect 170234 34226 175735 34288
rect 170873 33979 175639 34041
rect 176826 29656 187502 29718
rect 176826 29110 176910 29656
rect 187414 29110 187502 29656
rect 176826 29030 187502 29110
rect 175492 26516 176029 26596
rect 175492 24915 175555 26516
rect 175954 24915 176029 26516
rect 175492 24840 176029 24915
rect 176576 26528 177113 26591
rect 176576 24927 176639 26528
rect 177038 24927 177113 26528
rect 176576 24835 177113 24927
rect 137650 11398 137884 11418
rect 137650 10966 137668 11398
rect 137868 10966 137884 11398
rect 137650 10940 137884 10966
rect 137974 11396 138208 11418
rect 137974 10964 137992 11396
rect 138192 10964 138208 11396
rect 137974 10940 138208 10964
rect 166910 11412 167140 11430
rect 166910 10970 166932 11412
rect 167118 10970 167140 11412
rect 166910 10946 167140 10970
rect 167200 11410 167430 11432
rect 167200 10968 167222 11410
rect 167408 10968 167430 11410
rect 167200 10948 167430 10968
rect 136762 8396 190046 8406
rect 136762 8289 172516 8396
rect 172752 8289 190046 8396
rect 136762 8278 190046 8289
rect 136762 7932 190046 8132
rect 136762 7772 190046 7784
rect 136762 7665 172508 7772
rect 172744 7665 190046 7772
rect 136762 7656 190046 7665
rect 136762 7310 190046 7510
rect 136762 7151 190046 7162
rect 136762 7044 172508 7151
rect 172744 7044 190046 7151
rect 136762 7034 190046 7044
<< via3 >>
rect 153572 60458 155089 60810
rect 150103 59834 151655 60183
rect 181062 34968 187436 35554
rect 176910 29110 187414 29656
rect 175555 24915 175954 26516
rect 176639 24927 177038 26528
rect 137668 10966 137868 11398
rect 137992 10964 138192 11396
rect 166932 10970 167118 11412
rect 167222 10968 167408 11410
rect 148574 10488 149640 10809
rect 156116 9884 157197 10215
rect 172516 8289 172752 8396
rect 172508 7665 172744 7772
rect 172508 7044 172744 7151
<< metal4 >>
rect 192853 69022 193914 69106
rect 192853 67944 192943 69022
rect 193812 67944 193914 69022
rect 153550 64947 155115 65290
rect 153550 63632 153658 64947
rect 155009 63632 155115 64947
rect 150076 62801 151681 63222
rect 150076 61486 150206 62801
rect 151557 61486 151681 62801
rect 150076 60183 151681 61486
rect 153550 60810 155115 63632
rect 191197 64959 191960 65135
rect 191197 63620 191253 64959
rect 191878 63620 191960 64959
rect 153550 60458 153572 60810
rect 155089 60458 155115 60810
rect 153550 60423 155115 60458
rect 171674 62799 172694 63062
rect 171674 61472 171742 62799
rect 172605 61472 172694 62799
rect 150076 59834 150103 60183
rect 151655 59834 151681 60183
rect 150076 59795 151681 59834
rect 171674 35885 172694 61472
rect 171674 35554 187598 35885
rect 171674 34968 181062 35554
rect 187436 34968 187598 35554
rect 171674 34865 187598 34968
rect 137648 11398 137885 11418
rect 137648 10966 137668 11398
rect 137868 10966 137885 11398
rect 137648 8001 137885 10966
rect 137973 11396 138210 11416
rect 137973 10964 137992 11396
rect 138192 10964 138210 11396
rect 137973 7312 138210 10964
rect 166910 11412 167140 11430
rect 166910 10970 166932 11412
rect 167118 10970 167140 11412
rect 166910 10946 167140 10970
rect 167200 11410 167430 11432
rect 167200 10968 167222 11410
rect 167408 10968 167430 11410
rect 167200 10948 167430 10968
rect 148524 10809 149674 10843
rect 148524 10488 148574 10809
rect 149640 10488 149674 10809
rect 148524 2174 149674 10488
rect 156059 10215 157241 10309
rect 156059 9884 156116 10215
rect 157197 9884 157241 10215
rect 156059 9849 157241 9884
rect 156076 4568 157235 9849
rect 166912 7336 167138 10946
rect 167200 7953 167426 10948
rect 172498 8396 172765 34865
rect 191197 29792 191960 63620
rect 176805 29656 191960 29792
rect 176805 29110 176910 29656
rect 187414 29110 191960 29656
rect 176805 29029 191960 29110
rect 172498 8289 172516 8396
rect 172752 8289 172765 8396
rect 172498 7772 172765 8289
rect 172498 7665 172508 7772
rect 172744 7665 172765 7772
rect 172498 7151 172765 7665
rect 172498 7044 172508 7151
rect 172744 7044 172765 7151
rect 172498 7004 172765 7044
rect 175492 26516 176029 26596
rect 175492 24915 175555 26516
rect 175954 24915 176029 26516
rect 156076 3217 156181 4568
rect 157121 3217 157235 4568
rect 156076 3072 157235 3217
rect 148524 823 148622 2174
rect 149562 823 149674 2174
rect 148524 580 149674 823
rect 175492 2221 176029 24915
rect 176576 26528 177113 26591
rect 176576 24927 176639 26528
rect 177038 24927 177113 26528
rect 176576 4639 177113 24927
rect 176576 3211 176649 4639
rect 177032 3211 177113 4639
rect 176576 3132 177113 3211
rect 192853 4612 193914 67944
rect 192853 3207 192931 4612
rect 193816 3207 193914 4612
rect 192853 3072 193914 3207
rect 194710 67091 195771 67236
rect 194710 65970 194788 67091
rect 195667 65970 195771 67091
rect 175492 776 175531 2221
rect 175973 776 176029 2221
rect 175492 660 176029 776
rect 194710 2206 195771 65970
rect 194710 801 194793 2206
rect 195678 801 195771 2206
rect 194710 566 195771 801
<< via4 >>
rect 192943 67944 193812 69022
rect 153658 63632 155009 64947
rect 150206 61486 151557 62801
rect 191253 63620 191878 64959
rect 171742 61472 172605 62799
rect 156181 3217 157121 4568
rect 148622 823 149562 2174
rect 176649 3211 177032 4639
rect 192931 3207 193816 4612
rect 194788 65970 195667 67091
rect 175531 776 175973 2221
rect 194793 801 195678 2206
<< metal5 >>
rect 134778 69022 193994 69105
rect 134778 67944 192943 69022
rect 193812 67944 193994 69022
rect 134778 67852 193994 67944
rect 134816 67091 195923 67168
rect 134816 65970 194788 67091
rect 195667 65970 195923 67091
rect 134816 65915 195923 65970
rect 134593 64959 193084 65030
rect 134593 64947 191253 64959
rect 134593 63632 153658 64947
rect 155009 63632 191253 64947
rect 134593 63620 191253 63632
rect 191878 63620 193084 64959
rect 134593 63536 193084 63620
rect 134806 62801 193297 62895
rect 134806 61486 150206 62801
rect 151557 62799 193297 62801
rect 151557 61486 171742 62799
rect 134806 61472 171742 61486
rect 172605 61472 193297 62799
rect 134806 61401 193297 61472
rect 136826 4639 195936 4706
rect 136826 4568 176649 4639
rect 136826 3217 156181 4568
rect 157121 3217 176649 4568
rect 136826 3211 176649 3217
rect 177032 4612 195936 4639
rect 177032 3211 192931 4612
rect 136826 3207 192931 3211
rect 193816 3207 195936 4612
rect 136826 3138 195936 3207
rect 136826 2221 195980 2281
rect 136826 2174 175531 2221
rect 136826 823 148622 2174
rect 149562 823 175531 2174
rect 136826 776 175531 823
rect 175973 2206 195980 2221
rect 175973 801 194793 2206
rect 195678 801 195980 2206
rect 175973 776 195980 801
rect 136826 713 195980 776
use cv3_via2_8cut  cv3_via2_8cut_0
timestamp 1719106786
transform 1 0 168744 0 1 -28464
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_43
timestamp 1719106786
transform 1 0 168742 0 1 -27984
box 6850 62208 6998 62544
use cv3_via3_30cut  cv3_via3_30cut_181
timestamp 1719173267
transform 0 1 45904 -1 0 574842
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_182
timestamp 1719173267
transform 0 1 76043 -1 0 574838
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_183
timestamp 1719173267
transform 0 1 75669 -1 0 574209
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_184
timestamp 1719173267
transform 0 1 46273 -1 0 574213
box 566656 91154 566956 91980
use cv3_via_3cut  cv3_via_3cut_133
timestamp 1719452912
transform 1 0 165723 0 1 -105170
box 10601 106968 10663 107172
use sky130_ef_ip__cdac3v_12bit  sky130_ef_ip__cdac3v_12bit_0 ../ip/sky130_ef_ip__cdac3v_12bit/mag
timestamp 1731119720
transform 1 0 81345 0 -1 24388
box 52849 -36568 89580 15691
use sky130_ef_ip__scomp3v  sky130_ef_ip__scomp3v_0 ../ip/sky130_ef_ip__ccomp3v/mag
timestamp 1731119720
transform -1 0 187546 0 -1 32814
box -58 -3122 11186 4094
<< labels >>
flabel metal2 153040 0 153068 300 0 FreeSans 240 90 0 0 adc0_dac_val_11
port 640 nsew
flabel metal2 152928 0 152956 300 0 FreeSans 240 90 0 0 adc0_dac_val_10
port 641 nsew
flabel metal2 152816 0 152844 300 0 FreeSans 240 90 0 0 adc0_dac_val_9
port 642 nsew
flabel metal2 152704 0 152732 300 0 FreeSans 240 90 0 0 adc0_dac_val_8
port 643 nsew
flabel metal2 152592 0 152620 300 0 FreeSans 240 90 0 0 adc0_dac_val_7
port 644 nsew
flabel metal2 152480 0 152508 300 0 FreeSans 240 90 0 0 adc0_dac_val_6
port 645 nsew
flabel metal2 152368 0 152396 300 0 FreeSans 240 90 0 0 adc0_dac_val_5
port 646 nsew
flabel metal2 152256 0 152284 300 0 FreeSans 240 90 0 0 adc0_dac_val_4
port 647 nsew
flabel metal2 152144 0 152172 300 0 FreeSans 240 90 0 0 adc0_dac_val_3
port 648 nsew
flabel metal2 152032 0 152060 300 0 FreeSans 240 90 0 0 adc0_dac_val_2
port 649 nsew
flabel metal2 151920 0 151948 300 0 FreeSans 240 90 0 0 adc0_dac_val_1
port 650 nsew
flabel metal2 151808 0 151836 300 0 FreeSans 240 90 0 0 adc0_dac_val_0
port 651 nsew
flabel metal1 136762 8478 136866 8514 0 FreeSans 320 0 0 0 adc0_ena
port 652 nsew
flabel metal2 150226 102 150262 256 0 FreeSans 320 90 0 0 adc0_reset
port 653 nsew
flabel metal1 170288 1969 170425 2005 0 FreeSans 320 0 0 0 adc0_comp_out
port 654 nsew
flabel metal1 170288 1885 170426 1921 0 FreeSans 320 0 0 0 adc0_hold
port 656 nsew
flabel metal3 136762 7932 137018 8132 0 FreeSans 320 0 0 0 adc_vrefH
port 657 nsew
flabel metal3 136762 7310 137137 7510 0 FreeSans 320 0 0 0 adc_vrefL
port 658 nsew
flabel metal5 171792 3138 172938 4704 0 FreeSans 1600 0 0 0 vccd0
port 659 nsew
flabel metal5 171586 713 172629 2279 0 FreeSans 1600 0 0 0 vssd0
port 660 nsew
flabel metal5 134965 61518 136829 62782 0 FreeSans 1600 0 0 0 vssa0
port 663 nsew
flabel metal5 134751 63658 136615 64922 0 FreeSans 1600 0 0 0 vdda0
port 664 nsew
flabel metal3 174483 34002 174491 34011 0 FreeSans 800 0 0 0 adc_aval
<< end >>
